module top_module ( input a, input b, output out );
    
    mod_a instance1 ( a, b, out );

endmodule
